module btog(g,b);
input[3:0]b;
output[3:0]g;
 buf buf_g1(g[3],b[3]);
 xor xor_g1(g[2],b[3],b[2]);
 xor xor_g2(g[1],b[2],b[1]);
 xor xor_g3(g[0],b[1],b[0]);
endmodule
